* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT halfadder S X Y VDD GND C
** N=13 EP=6 IP=0 FDC=18
M0 6 Y GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=2605 $Y=775 $D=0
M1 S X 2 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=4620 $Y=255 $D=0
M2 2 6 S GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=5310 $Y=255 $D=0
M3 GND Y 2 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=6000 $Y=255 $D=0
M4 2 7 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=6690 $Y=255 $D=0
M5 GND X 7 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=8700 $Y=775 $D=0
M6 10 X 5 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=10710 $Y=840 $D=0
M7 GND Y 10 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=11400 $Y=840 $D=0
M8 C 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=13415 $Y=845 $D=0
M9 6 Y VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=2620 $Y=2275 $D=1
M10 12 X VDD VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=4.9e-13 PD=7.4e-07 PS=1.98e-06 $X=4630 $Y=2275 $D=1
M11 S 6 12 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.7e-13 PD=5.1e-07 PS=7.4e-07 $X=5550 $Y=2275 $D=1
M12 13 Y S VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=2.55e-13 PD=2.5e-07 PS=5.1e-07 $X=6240 $Y=2275 $D=1
M13 VDD 7 13 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.25e-13 PD=1.98e-06 PS=2.5e-07 $X=6670 $Y=2275 $D=1
M14 VDD X 7 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=8680 $Y=2275 $D=1
M15 5 X VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=10705 $Y=2275 $D=1
M16 VDD Y 5 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=11400 $Y=2275 $D=1
M17 C 5 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=13415 $Y=2275 $D=1
.ENDS
***************************************
