* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT fourbitsadder A0 B0 S0 C0 A1 B1 S1 A2 B2 S2 A3 B3 S3 GND VDD C4
** N=95 EP=16 IP=0 FDC=168
M0 49 B0 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=5415 $Y=7665 $D=0
M1 16 A0 8 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=6875 $Y=7665 $D=0
M2 8 49 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=7565 $Y=7665 $D=0
M3 GND B0 8 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8255 $Y=7665 $D=0
M4 8 50 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=8945 $Y=7665 $D=0
M5 GND A0 50 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=10955 $Y=8185 $D=0
M6 51 A0 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=12415 $Y=8185 $D=0
M7 11 B0 51 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=13105 $Y=8185 $D=0
M8 1 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=14570 $Y=8185 $D=0
M9 GND 12 17 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=16030 $Y=8185 $D=0
M10 52 16 12 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=17495 $Y=8185 $D=0
M11 GND C0 52 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=18185 $Y=8185 $D=0
M12 53 C0 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=19645 $Y=8185 $D=0
M13 GND 53 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=21655 $Y=7665 $D=0
M14 15 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=22345 $Y=7665 $D=0
M15 S0 54 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=23035 $Y=7665 $D=0
M16 15 C0 S0 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=23725 $Y=7665 $D=0
M17 GND 16 54 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=25185 $Y=7665 $D=0
M18 18 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=26645 $Y=7665 $D=0
M19 GND 1 18 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=27335 $Y=7665 $D=0
M20 2 18 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=28800 $Y=7665 $D=0
M21 56 B1 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=30260 $Y=7665 $D=0
M22 26 A1 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=31720 $Y=7665 $D=0
M23 19 56 26 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=32410 $Y=7665 $D=0
M24 GND B1 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=33100 $Y=7665 $D=0
M25 19 57 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=33790 $Y=7665 $D=0
M26 GND A1 57 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=35800 $Y=8185 $D=0
M27 58 A1 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=37260 $Y=8185 $D=0
M28 22 B1 58 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=37950 $Y=8185 $D=0
M29 3 22 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=39415 $Y=8185 $D=0
M30 GND 23 27 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=40875 $Y=8185 $D=0
M31 59 26 23 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=42340 $Y=8185 $D=0
M32 GND 2 59 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=43030 $Y=8185 $D=0
M33 60 2 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=44490 $Y=8185 $D=0
M34 GND 60 25 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=46500 $Y=7665 $D=0
M35 25 26 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=47190 $Y=7665 $D=0
M36 S1 61 25 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=47880 $Y=7665 $D=0
M37 25 2 S1 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=48570 $Y=7665 $D=0
M38 GND 26 61 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=50030 $Y=7665 $D=0
M39 28 27 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=51490 $Y=7665 $D=0
M40 GND 3 28 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=52180 $Y=7665 $D=0
M41 4 28 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=53645 $Y=7665 $D=0
M42 63 B2 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=55105 $Y=7665 $D=0
M43 36 A2 29 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=56565 $Y=7665 $D=0
M44 29 63 36 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=57255 $Y=7665 $D=0
M45 GND B2 29 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=57945 $Y=7665 $D=0
M46 29 64 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=58635 $Y=7665 $D=0
M47 GND A2 64 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=60645 $Y=8185 $D=0
M48 65 A2 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=62105 $Y=8185 $D=0
M49 32 B2 65 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=62795 $Y=8185 $D=0
M50 5 32 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=64260 $Y=8185 $D=0
M51 GND 33 37 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=65720 $Y=8185 $D=0
M52 66 36 33 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=67185 $Y=8185 $D=0
M53 GND 4 66 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=67875 $Y=8185 $D=0
M54 67 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=69335 $Y=8185 $D=0
M55 GND 67 35 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=71345 $Y=7665 $D=0
M56 35 36 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=72035 $Y=7665 $D=0
M57 S2 68 35 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=72725 $Y=7665 $D=0
M58 35 4 S2 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=73415 $Y=7665 $D=0
M59 GND 36 68 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=74875 $Y=7665 $D=0
M60 38 37 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=76335 $Y=7665 $D=0
M61 GND 5 38 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=77025 $Y=7665 $D=0
M62 6 38 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=78490 $Y=7665 $D=0
M63 70 B3 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=79950 $Y=7665 $D=0
M64 46 A3 39 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=81410 $Y=7665 $D=0
M65 39 70 46 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=82100 $Y=7665 $D=0
M66 GND B3 39 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=82790 $Y=7665 $D=0
M67 39 71 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=83480 $Y=7665 $D=0
M68 GND A3 71 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=85490 $Y=8185 $D=0
M69 72 A3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=86950 $Y=8185 $D=0
M70 42 B3 72 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=87640 $Y=8185 $D=0
M71 7 42 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=89105 $Y=8185 $D=0
M72 GND 43 47 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=90565 $Y=8185 $D=0
M73 73 46 43 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=92030 $Y=8185 $D=0
M74 GND 6 73 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=92720 $Y=8185 $D=0
M75 74 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=94180 $Y=8185 $D=0
M76 GND 74 45 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=96190 $Y=7665 $D=0
M77 45 46 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=96880 $Y=7665 $D=0
M78 S3 75 45 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=97570 $Y=7665 $D=0
M79 45 6 S3 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=98260 $Y=7665 $D=0
M80 GND 46 75 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=99720 $Y=7665 $D=0
M81 48 47 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=101180 $Y=7665 $D=0
M82 GND 7 48 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=101870 $Y=7665 $D=0
M83 C4 48 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=103335 $Y=7665 $D=0
M84 49 B0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=5425 $Y=9685 $D=1
M85 80 A0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=4.9e-13 PD=7.4e-07 PS=1.98e-06 $X=6885 $Y=9685 $D=1
M86 16 49 80 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.7e-13 PD=5.1e-07 PS=7.4e-07 $X=7805 $Y=9685 $D=1
M87 81 B0 16 VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=2.55e-13 PD=2.5e-07 PS=5.1e-07 $X=8495 $Y=9685 $D=1
M88 VDD 50 81 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.25e-13 PD=1.98e-06 PS=2.5e-07 $X=8925 $Y=9685 $D=1
M89 VDD A0 50 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=10935 $Y=9685 $D=1
M90 11 A0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=12395 $Y=9685 $D=1
M91 VDD B0 11 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=13090 $Y=9685 $D=1
M92 1 11 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=14550 $Y=9685 $D=1
M93 VDD 12 17 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=16050 $Y=9685 $D=1
M94 12 16 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=17510 $Y=9685 $D=1
M95 VDD C0 12 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=18205 $Y=9685 $D=1
M96 53 C0 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=19665 $Y=9685 $D=1
M97 82 53 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=4.9e-13 PD=2.5e-07 PS=1.98e-06 $X=21675 $Y=9685 $D=1
M98 S0 16 82 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=1.25e-13 PD=5.1e-07 PS=2.5e-07 $X=22105 $Y=9685 $D=1
M99 83 54 S0 VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=2.55e-13 PD=7.4e-07 PS=5.1e-07 $X=22795 $Y=9685 $D=1
M100 VDD C0 83 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.7e-13 PD=1.98e-06 PS=7.4e-07 $X=23715 $Y=9685 $D=1
M101 VDD 16 54 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=25175 $Y=9685 $D=1
M102 55 17 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=26645 $Y=9685 $D=1
M103 18 1 55 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=27340 $Y=9685 $D=1
M104 2 18 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=28800 $Y=9685 $D=1
M105 56 B1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=30270 $Y=9685 $D=1
M106 84 A1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=4.9e-13 PD=7.4e-07 PS=1.98e-06 $X=31730 $Y=9685 $D=1
M107 26 56 84 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.7e-13 PD=5.1e-07 PS=7.4e-07 $X=32650 $Y=9685 $D=1
M108 85 B1 26 VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=2.55e-13 PD=2.5e-07 PS=5.1e-07 $X=33340 $Y=9685 $D=1
M109 VDD 57 85 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.25e-13 PD=1.98e-06 PS=2.5e-07 $X=33770 $Y=9685 $D=1
M110 VDD A1 57 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=35780 $Y=9685 $D=1
M111 22 A1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=37240 $Y=9685 $D=1
M112 VDD B1 22 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=37935 $Y=9685 $D=1
M113 3 22 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=39395 $Y=9685 $D=1
M114 VDD 23 27 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=40895 $Y=9685 $D=1
M115 23 26 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=42355 $Y=9685 $D=1
M116 VDD 2 23 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=43050 $Y=9685 $D=1
M117 60 2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=44510 $Y=9685 $D=1
M118 86 60 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=4.9e-13 PD=2.5e-07 PS=1.98e-06 $X=46520 $Y=9685 $D=1
M119 S1 26 86 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=1.25e-13 PD=5.1e-07 PS=2.5e-07 $X=46950 $Y=9685 $D=1
M120 87 61 S1 VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=2.55e-13 PD=7.4e-07 PS=5.1e-07 $X=47640 $Y=9685 $D=1
M121 VDD 2 87 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.7e-13 PD=1.98e-06 PS=7.4e-07 $X=48560 $Y=9685 $D=1
M122 VDD 26 61 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=50020 $Y=9685 $D=1
M123 62 27 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=51490 $Y=9685 $D=1
M124 28 3 62 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=52185 $Y=9685 $D=1
M125 4 28 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=53645 $Y=9685 $D=1
M126 63 B2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=55115 $Y=9685 $D=1
M127 88 A2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=4.9e-13 PD=7.4e-07 PS=1.98e-06 $X=56575 $Y=9685 $D=1
M128 36 63 88 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.7e-13 PD=5.1e-07 PS=7.4e-07 $X=57495 $Y=9685 $D=1
M129 89 B2 36 VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=2.55e-13 PD=2.5e-07 PS=5.1e-07 $X=58185 $Y=9685 $D=1
M130 VDD 64 89 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.25e-13 PD=1.98e-06 PS=2.5e-07 $X=58615 $Y=9685 $D=1
M131 VDD A2 64 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=60625 $Y=9685 $D=1
M132 32 A2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=62085 $Y=9685 $D=1
M133 VDD B2 32 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=62780 $Y=9685 $D=1
M134 5 32 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=64240 $Y=9685 $D=1
M135 VDD 33 37 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=65740 $Y=9685 $D=1
M136 33 36 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=67200 $Y=9685 $D=1
M137 VDD 4 33 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=67895 $Y=9685 $D=1
M138 67 4 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=69355 $Y=9685 $D=1
M139 90 67 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=4.9e-13 PD=2.5e-07 PS=1.98e-06 $X=71365 $Y=9685 $D=1
M140 S2 36 90 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=1.25e-13 PD=5.1e-07 PS=2.5e-07 $X=71795 $Y=9685 $D=1
M141 91 68 S2 VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=2.55e-13 PD=7.4e-07 PS=5.1e-07 $X=72485 $Y=9685 $D=1
M142 VDD 4 91 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.7e-13 PD=1.98e-06 PS=7.4e-07 $X=73405 $Y=9685 $D=1
M143 VDD 36 68 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=74865 $Y=9685 $D=1
M144 69 37 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=76335 $Y=9685 $D=1
M145 38 5 69 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=77030 $Y=9685 $D=1
M146 6 38 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=78490 $Y=9685 $D=1
M147 70 B3 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=79960 $Y=9685 $D=1
M148 92 A3 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=4.9e-13 PD=7.4e-07 PS=1.98e-06 $X=81420 $Y=9685 $D=1
M149 46 70 92 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.7e-13 PD=5.1e-07 PS=7.4e-07 $X=82340 $Y=9685 $D=1
M150 93 B3 46 VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=2.55e-13 PD=2.5e-07 PS=5.1e-07 $X=83030 $Y=9685 $D=1
M151 VDD 71 93 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.25e-13 PD=1.98e-06 PS=2.5e-07 $X=83460 $Y=9685 $D=1
M152 VDD A3 71 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=85470 $Y=9685 $D=1
M153 42 A3 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=86930 $Y=9685 $D=1
M154 VDD B3 42 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=87625 $Y=9685 $D=1
M155 7 42 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=89085 $Y=9685 $D=1
M156 VDD 43 47 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=90585 $Y=9685 $D=1
M157 43 46 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=92045 $Y=9685 $D=1
M158 VDD 6 43 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=92740 $Y=9685 $D=1
M159 74 6 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=94200 $Y=9685 $D=1
M160 94 74 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=4.9e-13 PD=2.5e-07 PS=1.98e-06 $X=96210 $Y=9685 $D=1
M161 S3 46 94 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=1.25e-13 PD=5.1e-07 PS=2.5e-07 $X=96640 $Y=9685 $D=1
M162 95 75 S3 VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=2.55e-13 PD=7.4e-07 PS=5.1e-07 $X=97330 $Y=9685 $D=1
M163 VDD 6 95 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=3.7e-13 PD=1.98e-06 PS=7.4e-07 $X=98250 $Y=9685 $D=1
M164 VDD 46 75 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=99710 $Y=9685 $D=1
M165 76 47 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=101180 $Y=9685 $D=1
M166 48 7 76 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=101875 $Y=9685 $D=1
M167 C4 48 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=103335 $Y=9685 $D=1
.ENDS
***************************************
