* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT XOR Y X F VDD GND
** N=10 EP=5 IP=0 FDC=12
M0 4 Y GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=14005 $Y=5060 $D=0
M1 F X 5 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=16005 $Y=3830 $D=0
M2 5 4 F GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=16695 $Y=3830 $D=0
M3 GND Y 5 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=17385 $Y=3830 $D=0
M4 5 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=18075 $Y=3830 $D=0
M5 GND X 6 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=20065 $Y=5060 $D=0
M6 4 Y VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=14005 $Y=6560 $D=1
M7 9 X VDD VDD P_18 L=1.8e-07 W=1e-06 AD=3.7e-13 AS=4.9e-13 PD=7.4e-07 PS=1.98e-06 $X=16015 $Y=6560 $D=1
M8 F 4 9 VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=3.7e-13 PD=5.1e-07 PS=7.4e-07 $X=16935 $Y=6560 $D=1
M9 10 Y F VDD P_18 L=1.8e-07 W=1e-06 AD=1.25e-13 AS=2.55e-13 PD=2.5e-07 PS=5.1e-07 $X=17625 $Y=6560 $D=1
M10 VDD 6 10 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=1.25e-13 PD=1.98e-06 PS=2.5e-07 $X=18055 $Y=6560 $D=1
M11 VDD X 6 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06 $X=20065 $Y=6560 $D=1
.ENDS
***************************************
