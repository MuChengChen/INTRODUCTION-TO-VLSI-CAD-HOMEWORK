*inverter*
.subckt inv in out_1 VDD GND

MpMos out_1 in VDD VDD p_18 W=1u L=0.18u
MnMos out_1 in GND GND n_18 W=0.5u L=0.18u

.ends


*nand*
.subckt nand A B out_2 VDD GND
MpMos1 out_2 A VDD VDD p_18 W=1u L=0.18u
MpMos2 out_2 B VDD VDD p_18 W=1u L=0.18u
MnMos1 out_2 A nMos2_D GND n_18 W=0.5u L=0.18u
MnMos2 nMos2_D B GND GND n_18 W=0.5u L=0.18u

.ends


*nor*
.subckt nor C D out_3 VDD GND
MpMos3 pMos3_D C VDD VDD p_18 W=1u L=0.18u
MpMos4 out_3 D pMos3_D VDD p_18 W=1u L=0.18u
MnMos3 out_3 D GND GND n_18 W=0.5u L=0.18u
MnMos4 out_3 C GND GND n_18 W=0.5u L=0.18u


.ends
