* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT DFF clk reset QX Q GND VDD D
** N=21 EP=7 IP=0 FDC=32
M0 14 clk GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=11485 $Y=16935 $D=0
M1 15 6 14 GND N_18 L=1.8e-07 W=5e-07 AD=1.2875e-13 AS=1.275e-13 PD=5.15e-07 PS=5.1e-07 $X=12175 $Y=16935 $D=0
M2 4 1 15 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.2875e-13 PD=1.48e-06 PS=5.15e-07 $X=12870 $Y=16935 $D=0
M3 11 1 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=14880 $Y=16935 $D=0
M4 2 6 11 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=15570 $Y=16935 $D=0
M5 16 2 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=17585 $Y=16940 $D=0
M6 17 clk 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.2875e-13 AS=1.275e-13 PD=5.15e-07 PS=5.1e-07 $X=18275 $Y=16940 $D=0
M7 6 reset 17 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.2875e-13 PD=1.48e-06 PS=5.15e-07 $X=18970 $Y=16940 $D=0
M8 18 reset GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=20980 $Y=16940 $D=0
M9 19 D 18 GND N_18 L=1.8e-07 W=5e-07 AD=1.2875e-13 AS=1.275e-13 PD=5.15e-07 PS=5.1e-07 $X=21670 $Y=16940 $D=0
M10 1 4 19 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.2875e-13 PD=1.48e-06 PS=5.15e-07 $X=22365 $Y=16940 $D=0
M11 20 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=24375 $Y=16940 $D=0
M12 21 reset 20 GND N_18 L=1.8e-07 W=5e-07 AD=1.2875e-13 AS=1.275e-13 PD=5.15e-07 PS=5.1e-07 $X=25065 $Y=16940 $D=0
M13 QX Q 21 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.2875e-13 PD=1.48e-06 PS=5.15e-07 $X=25760 $Y=16940 $D=0
M14 13 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=27770 $Y=16935 $D=0
M15 Q QX 13 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=28460 $Y=16935 $D=0
M16 4 clk VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=11485 $Y=18370 $D=1
M17 VDD 6 4 VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=2.55e-13 PD=5.15e-07 PS=5.1e-07 $X=12175 $Y=18370 $D=1
M18 4 1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=12870 $Y=18370 $D=1
M19 2 1 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=14880 $Y=18370 $D=1
M20 VDD 6 2 VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=15575 $Y=18370 $D=1
M21 6 2 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=17585 $Y=18370 $D=1
M22 VDD clk 6 VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=2.55e-13 PD=5.15e-07 PS=5.1e-07 $X=18275 $Y=18370 $D=1
M23 6 reset VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=18970 $Y=18370 $D=1
M24 1 reset VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=20980 $Y=18370 $D=1
M25 VDD D 1 VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=2.55e-13 PD=5.15e-07 PS=5.1e-07 $X=21670 $Y=18370 $D=1
M26 1 4 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=22365 $Y=18370 $D=1
M27 QX 4 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06 $X=24375 $Y=18370 $D=1
M28 VDD reset QX VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=2.55e-13 PD=5.15e-07 PS=5.1e-07 $X=25065 $Y=18370 $D=1
M29 QX Q VDD VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=25760 $Y=18370 $D=1
M30 Q 6 VDD VDD P_18 L=1.8e-07 W=1e-06 AD=2.575e-13 AS=4.9e-13 PD=5.15e-07 PS=1.98e-06 $X=27770 $Y=18370 $D=1
M31 VDD QX Q VDD P_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.575e-13 PD=1.98e-06 PS=5.15e-07 $X=28465 $Y=18370 $D=1
.ENDS
***************************************
