*halfadder*
.subckt halfadder X Y S C VDD GND

MpMos1 X_inv X VDD VDD p_18 W=1u L=0.18u
MnMos1 X_inv X GND GND n_18 W=0.5u L=0.18u

MpMos2 Y_inv Y VDD VDD p_18 W=1u L=0.18u
MnMo2 Y_inv Y GND GND n_18 W=0.5u L=0.18u

MpMos3 VDD X pmos3 VDD p_18 W=1u L=0.18u
MpMos4 pmos3 Y_inv S VDD p_18 W=1u L=0.18u

MpMos5 VDD X_inv pmos5 VDD p_18 W=1u L=0.18u
MpMos6 pmos5 Y S VDD p_18 W=1u L=0.18u

MnMos3 S X nmos3 GND n_18 W=0.5u L=0.18u
MnMos4 nmos3 X_inv GND GND n_18 W=0.5u L=0.18u

MnMos5 S Y_inv nmos3 GND n_18 W=0.5u L=0.18u
MnMos6 nmos3 Y GND GND n_18 W=0.5u L=0.18u

MpMos7 C1 X VDD VDD p_18 W=1u L=0.18u
MpMos8 C1 Y VDD VDD p_18 W=1u L=0.18u
MnMos7 C1 X nMos2_D GND n_18 W=0.5u L=0.18u
MnMos8 nMos2_D Y GND GND n_18 W=0.5u L=0.18u

MpMos9 C C1 VDD VDD p_18 W=1u L=0.18u
MnMos9 C C1 GND GND n_18 W=0.5u L=0.18u

.ends
